
module residual
import types::*;
(
  input logic clk
 );
  endmodule : residual
