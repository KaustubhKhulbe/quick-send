package types;

    typedef enum logic [3:0] {
        READ,
        WRITE,
        IDLE
    } cpu_state_t;




endpackage




