module top_tb ();
    timeunit 1ps;
    timeprecision 1ps;
    wire dut;

    final begin
        $display("Monitor: Simulation finished");
    end

endmodule : top_tb
