module compress
(
 input logic clk,
 input logic rst,
 input types::residual_compress_reg cr_reg,
 output types::compress_commit_reg cc_reg
 );

  always_comb begin
    end

endmodule : compress
